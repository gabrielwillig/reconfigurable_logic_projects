-- Library IEEE;
-- use IEEE.std_logic_1164.all;
-- use IEEE.numeric_std.all;
-- -- Gabriel Freitas Willig
-- Entity digital_cronometer_tb is
-- end;
-- Architecture test of digital_cronometer_tb is
-- component digital_cronometer is
-- 	port(   
-- 		CLK              :   IN  std_logic;
-- 		SW_1             :   IN std_logic;
-- 		SW_2             :   IN std_logic;
-- 		SWITCH           :	 IN std_logic;
-- 		Q_M, Q_L         :   OUT std_logic_vector(3 downto 0);
-- 		Q_CENT_M, Q_CENT_L : OUT std_logic_vector(3 downto 0)
--     );
-- End component;
-- signal   RST:	        std_logic := '1';
-- signal   CLOCK:      		std_logic;
-- signal   SW1, SW2:   	std_logic := '0';
-- signal   M_SEC,L_SEC:	std_logic_vector(3 downto 0);
-- signal   M_CENT,L_CENT:	std_logic_vector(3 downto 0);

-- Begin
--     DUT: digital_cronometer port map(
--         CLK => CLOCK,
--         SW_1 => SW1,
--         SW_2 => SW2,
--         SWITCH => RST,
--         Q_M => M_SEC,
--         Q_L => L_SEC,
--         Q_CENT_M => M_CENT,
--         Q_CENT_L => L_CENT
--     );

--     Process
--     Begin
--         SW1 <= '1';
--         wait for 100 ns;
--         SW1 <= '0';
--         wait for 15 ns;
--         SW1 <= '1';
--         wait;
--         --wait for 10 ns;
-- 		    --SW2 <= '1';
-- 		    --wait for 20 ns;
-- 		    --SW2 <= '0';
-- 		    --wait for 20 ns;
--         --SW1 <= '0';
--         --wait;
--     End process;

--     process
--     begin
--       RST <= '1';
--       wait for 25 ns;
--       RST <= '0';
--       wait;
--     end process;

--     process
--     begin
--       while true loop
--         CLOCK <= '0';
--         wait for 10 ns;
--         CLOCK <= '1';
--         wait for 10 ns;
--       end loop;
--       wait;
--     end process;

-- end architecture;